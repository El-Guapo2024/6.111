module  pwm(
            input wire clk_in,
            input wire rst_in,
            input wire signed [7:0] level_in,
            input wire direction,
            output logic pwm_out
  );
 
endmodule
`default_nettype wire